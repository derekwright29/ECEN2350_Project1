module AND_D(x,y,out,en);
   input [3:0] x,y;
   output [3:0] out;
	input en;

	assign out = x & y;
	
endmodule // AND_D

module OR_D(x,y,out,en);
   input [3:0] x,y;
   output [3:0] out;
	input en;

	assign out = x | y;

endmodule // OR_D

module XOR_D(x,y,out,en);
   input [3:0] x,y;
   output [3:0] out;
	input en;

	assign out = x ^ y;
	
endmodule // XOR_D

module NOT_D(z,out,en);
   input [7:0] z;
   output [7:0] out;
	input en;

	assign out = ~z;
 
endmodule // NOT_D


   
